module main(input in, clk, clear, output out);
    reg [2:0]q;
    always_ff@(posedge clk or posedge clear)
        begin
            if(clear)
                q<=0;
            else
                begin
                if(q==0 && in==0)
                    q<=0;
                else if(q==0 && in==1)
                    q<=1;
                else
                if(q==1 && in==0)
                    q<=2;
                else if(q==1 && in==1)
                    q<=1;
                else
                if(q==2 && in==0)
                    q<=3;
                else if(q==2 && in==1)
                    q<=1;
                 else
                if(q==3 && in==0)
                    q<=0;
                else if(q==3 && in==1)
                    q<=4;
                else
                if(q==4 && in==0)
                    q<=0;
                else if(q==4 && in==1)
                    q<=1;
                end
         
        end  
    assign out = (q==4); 


endmodule


module tb;
    reg clk, clear, x;
    wire out;

    main uut(x,clk,clear,out);

    always #2 clk=~clk;

   initial begin
        $monitor("time=%0t,clk=%b, x=%b, clear=%b, out=%b",$time,clk, x,clear, out);
        clk=0;
        clear=1;
        x=0;
        #2 clear = 0;
        #4 x=1; //5
        #4 x=0; //9
        #4 x=0; //13
        #4 x=1; //17
        #4 x=0; //21
        #4 x=0; 
        #4 x=1; 
        #4 x=1; 
        #4 x=0; 
        #4 x=0; 
        #4 x=1;        
        #2$finish;
    end 

endmodule
